garofalo@larain1.ee.ethz.ch.125393:1544107630